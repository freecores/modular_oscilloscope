-- epp.vhd

	