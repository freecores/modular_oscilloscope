-- epp.vhd