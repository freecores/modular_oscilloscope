-- epp.vhd
-- M�dulo principal integrador
-- Peque�a modificaci�n de prueba