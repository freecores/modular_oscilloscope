-- ctrl.vhd